CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
110 0 30 100 9
0 71 1363 720
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1363 720
177209362 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 1002 476 0 1 11
0 5
0
0 0 21360 270
2 0V
-1 -19 13 -11
2 T3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 1606 374 0 1 11
0 23
0
0 0 21360 270
2 0V
-1 -19 13 -11
2 T2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 945 174 0 1 11
0 15
0
0 0 21360 270
2 0V
-1 -19 13 -11
2 T1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 624 79 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 782
2 5V
-6 -21 8 -13
1 S
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
9 Inverter~
13 877 508 0 2 22
0 5 6
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 NOT2
12 -4 40 4
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 3 0
1 U
5394 0 0
0
0
9 2-In AND~
219 913 450 0 3 22
0 6 7 4
0
0 0 624 692
6 74LS08
-21 -24 21 -16
4 AND6
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 6 0
1 U
7734 0 0
0
0
13 SR Flip-Flop~
219 679 572 0 4 9
0 5 3 9 7
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
7 timer1a
-24 -55 25 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
9914 0 0
0
0
7 Ground~
168 809 524 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
4 LED~
171 805 492 0 2 2
10 10 2
0
0 0 880 512
4 LED1
16 0 44 8
2 R3
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3549 0 0
0
0
9 2-In AND~
219 729 445 0 3 22
0 9 8 10
0
0 0 624 692
6 74LS08
-21 -24 21 -16
4 AND5
-18 -25 10 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 6 0
1 U
7931 0 0
0
0
9 2-In AND~
219 686 221 0 3 22
0 12 13 11
0
0 0 624 692
6 74LS08
-21 -24 21 -16
4 AND4
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 5 0
1 U
9325 0 0
0
0
7 Ground~
168 524 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
4 LED~
171 529 385 0 2 2
10 8 2
0
0 0 880 0
4 LED2
17 0 45 8
4 D180
17 -10 45 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3834 0 0
0
0
7 Ground~
168 531 94 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
4 LED~
171 529 155 0 2 2
10 13 2
0
0 0 880 180
4 LED2
16 0 44 8
2 D0
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7668 0 0
0
0
9 2-In AND~
219 785 169 0 3 22
0 11 18 14
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 AND2
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 251535339
65 0 0 0 4 4 2 0
1 U
4718 0 0
0
0
8 2-In OR~
219 329 216 0 3 22
0 4 22 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 OR6
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 251535339
65 0 0 0 4 1 4 0
1 U
3874 0 0
0
0
9 2-In AND~
219 428 282 0 3 22
0 19 3 22
0
0 0 624 512
6 74LS08
-21 -24 21 -16
4 AND1
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
6671 0 0
0
0
9 2-In AND~
219 880 118 0 3 22
0 17 16 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 AND3
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3789 0 0
0
0
9 Inverter~
13 855 195 0 2 22
0 15 16
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 NOT1
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 3 0
1 U
4871 0 0
0
0
13 SR Flip-Flop~
219 711 140 0 4 9
0 15 19 18 17
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
7 timer1a
-24 -55 25 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3750 0 0
0
0
7 Ground~
168 776 11 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8778 0 0
0
0
4 LED~
171 744 41 0 2 2
10 14 2
0
0 0 880 180
4 LED1
16 0 44 8
2 R1
23 -10 37 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
538 0 0
0
0
13 SR Flip-Flop~
219 429 378 0 4 9
0 20 4 3 8
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
4 F180
-14 -55 14 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
6843 0 0
0
0
13 SR Flip-Flop~
219 429 248 0 4 9
0 21 20 19 13
0
0 0 4720 0
4 SRFF
-14 -53 14 -45
2 F0
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3136 0 0
0
0
32
0 2 3 0 0 4224 0 0 7 18 0 3
469 360
469 554
655 554
2 0 4 0 0 4096 0 24 0 0 3 2
405 360
278 360
3 1 4 0 0 12416 0 6 17 0 0 6
934 450
1058 450
1058 629
278 629
278 207
316 207
1 0 5 0 0 12416 0 7 0 0 5 5
655 536
600 536
600 583
953 583
953 546
1 1 5 0 0 0 0 1 5 0 0 4
1002 488
1002 546
880 546
880 526
2 1 6 0 0 4224 0 5 6 0 0 3
880 490
880 459
889 459
4 2 7 0 0 12416 0 7 6 0 0 4
703 536
768 536
768 441
889 441
0 2 8 0 0 4224 0 0 10 20 0 4
529 341
694 341
694 436
705 436
3 1 9 0 0 8320 0 7 10 0 0 6
709 554
729 554
729 474
688 474
688 454
705 454
1 3 10 0 0 8320 0 9 10 0 0 3
809 482
809 445
750 445
1 2 2 0 0 4096 0 8 9 0 0 2
809 518
809 502
3 1 11 0 0 4224 0 11 16 0 0 4
707 221
812 221
812 178
803 178
1 1 12 0 0 4224 0 4 11 0 0 3
624 91
624 230
662 230
2 0 13 0 0 4224 0 11 0 0 15 2
662 212
531 212
1 4 13 0 0 128 0 15 25 0 0 3
531 165
531 212
453 212
2 1 2 0 0 8192 0 23 22 0 0 3
746 31
746 5
776 5
3 1 14 0 0 4224 0 16 23 0 0 7
758 169
758 63
747 63
747 56
741 56
741 51
746 51
3 2 3 0 0 128 0 24 18 0 0 4
459 360
469 360
469 291
448 291
2 1 2 0 0 4096 0 13 12 0 0 4
529 395
529 428
524 428
524 435
4 1 8 0 0 128 0 24 13 0 0 4
453 342
453 341
529 341
529 375
1 0 15 0 0 12416 0 21 0 0 23 6
687 104
666 104
666 75
975 75
975 207
945 207
2 2 16 0 0 8320 0 20 19 0 0 3
858 177
856 177
856 127
1 1 15 0 0 0 0 3 20 0 0 4
945 186
945 219
858 219
858 213
4 1 17 0 0 4224 0 21 19 0 0 4
735 104
850 104
850 109
856 109
2 3 18 0 0 12416 0 16 21 0 0 4
803 160
816 160
816 122
741 122
0 2 19 0 0 8320 0 0 21 32 0 4
459 249
585 249
585 122
687 122
2 1 2 0 0 4224 0 15 14 0 0 2
531 145
531 102
1 0 20 0 0 4096 0 24 0 0 29 2
405 342
372 342
3 2 20 0 0 12416 0 19 25 0 0 6
901 118
902 118
902 410
372 410
372 230
405 230
3 1 21 0 0 4224 0 17 25 0 0 4
362 216
399 216
399 212
405 212
3 2 22 0 0 4224 0 18 17 0 0 4
403 282
294 282
294 225
316 225
3 1 19 0 0 0 0 25 18 0 0 3
459 230
459 273
448 273
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
497 290 633 334
507 298 635 330
23 Acionando motor 
180�
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
339 101 491 125
349 109 493 125
18 Acionando motor 0�
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
966 398 1118 442
976 406 1120 438
23 Sa�da do timer de 
3s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
730 537 898 581
740 545 900 577
25 Entrada do timer de 
3s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
970 152 1138 176
980 160 1140 176
20 Sa�da do timer de 1s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
783 1 967 45
793 9 969 41
22 Entrada do timer de 1s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
608 24 664 48
618 32 666 48
6 Sensor
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2557198 1079360 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 5
0
263664 8550464 100 100 0 0
77 66 1307 246
0 395 1366 719
1307 66
77 66
1307 66
1307 246
0 0
4.53041e-315 0 4.95446e-315 4.95446e-315 4.53041e-315 4.53041e-315
12401 0
4 1e-006 5
1
676 271
0 11 0 0 1	0 33 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
